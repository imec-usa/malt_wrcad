* HNL Generated netlist of AA_fluxshut_top
* GLOBAL Parameters
.param amplitude = 0.700 frequency = 10G m_in = 0.1p
* GLOBAL Scaling Parameters
*.param Xac=1.0
*.param Xlcomp=1.0
*.param Xjcomp=1.0
.param Xl=1.0
.param Xj=1.0
*.param Xpdc=1.0
.param Xa=1.0
.param Xr=1.0
* Timing corner definitions
.param timingX = 1.0
.global 0
* Include Statements
.include my_models_spice.mod
*Subcircuits
.subckt aa_fluxshut a i0 i1 q
XL0 a i0 rql_inductor_scale l=7.4e-12
Loff i0 i1 'm_in'
XL2 i1 net04 rql_inductor_scale l=1.47e-11
XL1 net04 q rql_inductor_scale l=7.4e-12
Xb0 i0 net023 rql_rsj_scale jjmod=rql25 ic=0.07 icrn=1
Xb1 net04 net08 rql_rsj_scale jjmod=rql25 ic=0.07 icrn=1
Lg0 net023 0 1e-12
Lg1 net08 0 1e-12
.ends aa_fluxshut
.subckt g_terminate i ic1=0.050
XR0 i 0 rql_resistor_scale r='0.7/ic1'
.ends g_terminate
*Input stage
L1 na 0 'm_in'
XL0 net017 na rql_inductor_scale l='1e-12*l0'
Xb0 net015 net017 rql_rsj_scale jjmod=rql25 ic='b0' icrn=1
*Flux shuttle stages
XI1 net015 i1a i1b net06 aa_fluxshut
XI2 net06 i2a i2b net07 aa_fluxshut
XI3 net07 i3a i3b net08 aa_fluxshut
XI4 net08 i4a i4b net05 aa_fluxshut
XI5 net05 i5a i5b net09 aa_fluxshut
XI6 net09 i6a i6b net010 aa_fluxshut
XI7 net010 i7a i7b net03 aa_fluxshut
XI8 net03 i8a i8b net029 aa_fluxshut
XI9 net029 i9a i9b net018 aa_fluxshut
XI10 net018 i10a i10b net025 aa_fluxshut
XI11 net025 i11a i11b net020 aa_fluxshut
XI12 net020 i12a i12b net02 aa_fluxshut
*flux shuttle terminationXb1 net02 net04 rql_rsj_scale jjmod=rql25 ic='b1' icrn=1
Lg1 net04 0 1e-12
XI13 net02 g_terminate ic1=0.07
*output amp
XL2 net031 net030 rql_inductor_scale l=1e-12
XL3 net032 0 rql_inductor_scale l=1e-12
XL4 net029 net026 rql_inductor_scale l='1e-12*l45'
XL5 net024 net025 rql_inductor_scale l='1e-12*l45'
XL6 net030 oo rql_inductor_scale l=4e-10
XR0 net030 oo rql_resistor_scale r=50
Xb2 net030 net032 rql_rsj_scale jjmod=rql25 ic='b2' \
icrn='1.0*b2*0.07/(b2*0.07+b34*0.040)'
Xb3 net026 net031 phib3 rql_junction_scale area='b34' jjmod=rql25
Xb4 net024 net031 phib4 rql_junction_scale area='b34' jjmod=rql25
*Input source
Ia 0 na 'phi0/m_in*inoff' +\
pulse(0 'phi0/m_in*inipp' 170ps 20ps 20ps 80ps 1) +\
pulse(0 'phi0/m_in*inipp' 370ps 20ps 20ps 80ps 1) +\
pulse(0 'phi0/m_in*inipp' 570ps 20ps 20ps 80ps 1) +\
0
*Four phase clock sources
I1 i1a i1b sin(0 'phi0/m_in*Xac*amplitude' 10GHz 00ps)
I2 i2a i2b sin(0 'phi0/m_in*Xac*amplitude' 10GHz 25ps)
I3 i3a i3b sin(0 'phi0/m_in*Xac*amplitude' 10GHz 50ps)
I4 i4a i4b sin(0 'phi0/m_in*Xac*amplitude' 10GHz 75ps)
I5 i5a i5b sin(0 'phi0/m_in*Xac*amplitude' 10GHz 00ps)
I6 i6a i6b sin(0 'phi0/m_in*Xac*amplitude' 10GHz 25ps)
I7 i7a i7b sin(0 'phi0/m_in*Xac*amplitude' 10GHz 50ps)
I8 i8a i8b sin(0 'phi0/m_in*Xac*amplitude' 10GHz 75ps)
I9 i9a i9b sin(0 'phi0/m_in*Xac*amplitude' 10GHz 00ps)
I10 i10a i10b sin(0 'phi0/m_in*Xac*amplitude' 10GHz 25ps)
I11 i11a i11b sin(0 'phi0/m_in*Xac*amplitude' 10GHz 50ps)
I12 i12a i12b sin(0 'phi0/m_in*Xac*amplitude' 10GHz 75ps)
*Output source
Iout 0 oo pwl(0 0 20ps 'Xpdc*80uA')
Rout 0 oo 50
*Analysis definition
.tran 1ps 1000ps 0ps uic
.end
